----*-vhdl-*--------------------------------------------------------------------
-- PLOMB
-- Banc mémoire RAM générique à simple accès
--------------------------------------------------------------------------------
-- DO 4/2015
--------------------------------------------------------------------------------
-- 32 bits
--------------------------------------------------------------------------------

--##############################################################################
--## This source file is copyrighted. Read the "lic.txt" file before use.     ##
--## Experimental version. No warranty of any sort. All rights reserved.      ##
--##############################################################################

-- Initialisation Bootloader
-- VAR=5  : Bootloader SparcsStation5     : 4ko
-- VAR=20 : Bootloader SparcsStation10/20 : 4ko

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
use std.textio.all;

LIBRARY work;
USE work.base_pack.ALL;
USE work.plomb_pack.ALL;

--##############################################################################

ENTITY iram_ts IS
  GENERIC (
    VAR : natural := 1);
  PORT (
    mem_w : IN  type_pvc_w;
    mem_r : OUT type_pvc_r;
    
    -- Global
    clk      : IN std_logic;
    reset_n  : IN std_logic
    );
END ENTITY iram_ts;

ARCHITECTURE ts OF iram_ts IS

--------------------------------------------------------------------------------

  CONSTANT SIZE : natural := 2 ** 10;
  TYPE type_mem IS ARRAY(0 TO SIZE-1) OF uv8;

-- INSERTCONST
  CONSTANT INIT5_0 : type_mem:=(
    x"03",x"81",x"01",x"FF",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"27",x"81",x"A1",x"01",
    x"27",x"81",x"A1",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"01",x"01",x"81",x"81",x"01",x"01",x"81",x"81",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"03",x"82",x"81",x"81",x"03",x"81",x"03",x"84",
    x"C2",x"82",x"84",x"C2",x"82",x"84",x"C2",x"01",
    x"01",x"01",x"03",x"82",x"9C",x"BC",x"A0",x"E0",
    x"C1",x"05",x"84",x"07",x"86",x"82",x"01",x"40",
    x"01",x"01",x"03",x"84",x"C4",x"82",x"C2",x"01",
    x"01",x"81",x"01",x"03",x"81",x"03",x"81",x"01",
    x"A6",x"83",x"A1",x"82",x"81",x"81",x"01",x"01",
    x"01",x"E0",x"E4",x"E8",x"EC",x"F0",x"F4",x"F8",
    x"FC",x"81",x"82",x"81",x"81",x"01",x"01",x"01",
    x"A7",x"A1",x"A0",x"81",x"01",x"01",x"01",x"81",
    x"81",x"E0",x"E4",x"E8",x"EC",x"F0",x"F4",x"F8",
    x"FC",x"81",x"81",x"81",x"81",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"F0",x"02",x"01",x"07",
    x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"07",
    x"04",x"0B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
    x"D2",x"81",x"01",x"D2",x"81",x"01",x"D2",x"81",
    x"01",x"D0",x"81",x"01",x"D0",x"81",x"01",x"D0",
    x"81",x"01",x"03",x"82",x"C4",x"80",x"02",x"01",
    x"03",x"82",x"D0",x"81",x"01",x"03",x"84",x"10",
    x"82",x"C8",x"80",x"02",x"01",x"C6",x"90",x"C6",
    x"80",x"12",x"C6",x"81",x"01",x"03",x"82",x"C4",
    x"80",x"02",x"01",x"03",x"82",x"D0",x"81",x"01",
    x"84",x"03",x"82",x"C4",x"84",x"C4",x"84",x"C4",
    x"84",x"C4",x"86",x"C6",x"C0",x"C4",x"84",x"C4",
    x"C4",x"84",x"C4",x"84",x"C4",x"84",x"C4",x"81",
    x"01",x"03",x"82",x"C4",x"80",x"02",x"01",x"03",
    x"82",x"C2",x"80",x"08",x"84",x"84",x"03",x"85",
    x"82",x"C6",x"80",x"02",x"01",x"03",x"82",x"C2",
    x"90",x"80",x"18",x"90",x"82",x"90",x"81",x"01",
    x"9D",x"05",x"07",x"88",x"86",x"82",x"84",x"9B",
    x"DA",x"D8",x"80",x"02",x"01",x"DA",x"82",x"80",
    x"12",x"B1",x"81",x"81",x"03",x"C0",x"05",x"86",
    x"C6",x"C0",x"86",x"C6",x"C0",x"86",x"C6",x"C0",
    x"D2",x"88",x"C6",x"C0",x"80",x"02",x"07",x"C0",
    x"82",x"C2",x"C0",x"88",x"C8",x"C0",x"C2",x"C0",
    x"81",x"01",x"9D",x"03",x"88",x"C8",x"05",x"C0",
    x"86",x"C6",x"C0",x"9A",x"DA",x"C0",x"9A",x"DA",
    x"C0",x"C6",x"C0",x"C8",x"C0",x"C6",x"81",x"81",
    x"9D",x"03",x"84",x"C4",x"05",x"C0",x"86",x"C6",
    x"C0",x"86",x"C6",x"C0",x"86",x"C6",x"C0",x"C6",
    x"07",x"88",x"98",x"9A",x"86",x"D6",x"C0",x"D4",
    x"80",x"02",x"01",x"DA",x"80",x"02",x"01",x"C4",
    x"80",x"02",x"05",x"C0",x"86",x"C6",x"C0",x"88",
    x"C8",x"C0",x"C6",x"C0",x"81",x"81",x"9D",x"05",
    x"86",x"82",x"C6",x"86",x"C6",x"86",x"C6",x"86",
    x"C6",x"88",x"C8",x"C0",x"C6",x"86",x"C6",x"C6",
    x"86",x"C6",x"86",x"C6",x"88",x"86",x"84",x"C6",
    x"03",x"10",x"82",x"DA",x"80",x"02",x"01",x"C6",
    x"82",x"C6",x"80",x"12",x"C6",x"03",x"86",x"05",
    x"C6",x"82",x"80",x"12",x"01",x"05",x"03",x"86",
    x"82",x"10",x"84",x"DA",x"80",x"02",x"01",x"C8",
    x"82",x"C8",x"80",x"12",x"C8",x"23",x"35",x"37",
    x"39",x"3B",x"2F",x"2D",x"2B",x"B4",x"B6",x"B8",
    x"BA",x"AE",x"AC",x"AA",x"A4",x"A0",x"A8",x"C2",
    x"80",x"02",x"01",x"C2",x"82",x"80",x"12",x"80",
    x"05",x"03",x"86",x"82",x"10",x"84",x"DA",x"80",
    x"02",x"01",x"C8",x"82",x"C8",x"80",x"12",x"C8",
    x"81",x"81",x"12",x"80",x"82",x"07",x"05",x"C8",
    x"80",x"22",x"82",x"84",x"86",x"89",x"C8",x"DA",
    x"80",x"02",x"01",x"C8",x"84",x"80",x"32",x"83",
    x"82",x"10",x"84",x"C8",x"80",x"02",x"01",x"C6",
    x"82",x"C6",x"80",x"12",x"C6",x"03",x"84",x"10",
    x"82",x"80",x"12",x"01",x"03",x"84",x"10",x"82",
    x"C8",x"80",x"02",x"01",x"C6",x"82",x"C6",x"80",
    x"12",x"C6",x"82",x"10",x"84",x"C8",x"80",x"02",
    x"01",x"C6",x"82",x"C6",x"80",x"12",x"C6",x"A6",
    x"31",x"33",x"7F",x"90",x"7F",x"90",x"A6",x"80",
    x"12",x"82",x"10",x"84",x"C8",x"80",x"02",x"01",
    x"C6",x"82",x"C6",x"80",x"12",x"C6",x"A6",x"31",
    x"33",x"7F",x"90",x"A6",x"80",x"12",x"01",x"A6",
    x"B0",x"10",x"33",x"D2",x"90",x"93",x"A6",x"7F",
    x"93",x"80",x"0A",x"82",x"10",x"84",x"C8",x"80",
    x"02",x"01",x"C6",x"82",x"C6",x"80",x"12",x"C6",
    x"82",x"09",x"07",x"05",x"DA",x"D8",x"9B",x"99",
    x"80",x"22",x"82",x"84",x"86",x"89",x"C8",x"DA",
    x"80",x"02",x"01",x"C8",x"84",x"80",x"32",x"83",
    x"82",x"10",x"84",x"C8",x"80",x"02",x"01",x"C6",
    x"82",x"C6",x"80",x"12",x"C6",x"03",x"84",x"10",
    x"82",x"80",x"12",x"01",x"82",x"10",x"84",x"C8",
    x"80",x"02",x"01",x"C6",x"82",x"C6",x"80",x"12",
    x"C6",x"30",x"C8",x"80",x"02",x"01",x"C6",x"82",
    x"C6",x"80",x"12",x"C6",x"30",x"84",x"12",x"82",
    x"30",x"C8",x"80",x"02",x"01",x"C6",x"82",x"C6",
    x"80",x"12",x"C6",x"30",x"C2",x"80",x"02",x"03",
    x"82",x"C2",x"82",x"82",x"80",x"18",x"83",x"C2",
    x"81",x"01",x"C2",x"80",x"02",x"01",x"C2",x"80",
    x"02",x"80",x"12",x"01",x"30",x"C2",x"80",x"02",
    x"01",x"C2",x"80",x"02",x"80",x"12",x"01",x"30",
    x"7F",x"27",x"7F",x"B0",x"B0",x"F0",x"B2",x"7F",
    x"B0",x"B1",x"90",x"B0",x"10",x"A6",x"7F",x"B2",
    x"D0",x"A6",x"C2",x"80",x"0A",x"01",x"10",x"B0",
    x"7F",x"01",x"7F",x"B2",x"90",x"7F",x"A7",x"B2",
    x"B0",x"7F",x"F2",x"B0",x"90",x"B1",x"03",x"B0",
    x"27",x"B0",x"B2",x"10",x"A6",x"7F",x"B2",x"D0",
    x"A6",x"C2",x"80",x"0A",x"01",x"10",x"B0",x"7F",
    x"01",x"7F",x"B2",x"7F",x"A6",x"90",x"A7",x"7F",
    x"A6",x"A7",x"B2",x"B0",x"7F",x"F2",x"B0",x"90",
    x"B1",x"03",x"B0",x"27",x"B0",x"B2",x"10",x"A6",
    x"7F",x"B2",x"D0",x"A6",x"C2",x"80",x"0A",x"01",
    x"B0",x"80",x"2A",x"A4",x"7F",x"01",x"30",x"00",
    x"42",x"6C",x"65",x"00",x"3E",x"00",x"45",x"20",
    x"0A",x"00",x"0A",x"00",x"4E",x"42",x"4B",x"45",
    x"45",x"00",x"42",x"4B",x"46",x"48",x"49",x"0D",
    x"46",x"48",x"53",x"00",x"54",x"20",x"4F",x"00",
    x"54",x"20",x"0D",x"00",x"3E",x"00",x"30",x"34",
    x"38",x"43",x"00",x"30",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );

  CONSTANT INIT5_1 : type_mem:=(
    x"3C",x"C0",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"3C",x"C4",x"50",x"00",
    x"3C",x"C4",x"50",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"00",x"10",x"20",x"30",x"40",x"50",x"60",x"70",
    x"80",x"90",x"A0",x"B0",x"C0",x"D0",x"E0",x"F0",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"00",x"00",x"C4",x"CC",x"00",x"00",x"C4",x"CC",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"00",x"10",x"88",x"90",x"3C",x"98",x"3F",x"10",
    x"A0",x"10",x"10",x"A0",x"10",x"10",x"A0",x"00",
    x"00",x"00",x"3C",x"10",x"10",x"10",x"10",x"23",
    x"0B",x"3C",x"10",x"3C",x"10",x"10",x"00",x"00",
    x"00",x"00",x"3C",x"10",x"20",x"10",x"A0",x"00",
    x"00",x"C0",x"00",x"3C",x"98",x"00",x"C0",x"00",
    x"10",x"34",x"2C",x"14",x"E0",x"90",x"00",x"00",
    x"00",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",
    x"3B",x"E8",x"10",x"C4",x"CC",x"00",x"00",x"00",
    x"2C",x"34",x"14",x"94",x"00",x"00",x"00",x"E8",
    x"E8",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",
    x"1B",x"E0",x"E0",x"C4",x"CC",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"00",x"00",x"00",x"80",
    x"00",x"10",x"20",x"30",x"40",x"50",x"60",x"70",
    x"00",x"00",x"A0",x"B0",x"C0",x"D0",x"E0",x"F0",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"2A",x"C3",x"00",x"32",x"C3",x"00",x"22",x"C3",
    x"00",x"0A",x"C3",x"00",x"12",x"C3",x"00",x"02",
    x"C3",x"00",x"3C",x"10",x"08",x"88",x"BF",x"00",
    x"3C",x"10",x"28",x"C3",x"00",x"3C",x"10",x"80",
    x"10",x"08",x"89",x"BF",x"00",x"28",x"02",x"4A",
    x"A0",x"BF",x"0A",x"C3",x"00",x"3C",x"10",x"08",
    x"88",x"BF",x"00",x"3C",x"10",x"08",x"C3",x"00",
    x"10",x"3C",x"10",x"28",x"10",x"28",x"10",x"28",
    x"10",x"28",x"10",x"28",x"28",x"28",x"10",x"28",
    x"28",x"10",x"28",x"10",x"28",x"10",x"28",x"C3",
    x"00",x"3C",x"10",x"08",x"88",x"BF",x"00",x"3C",
    x"10",x"08",x"A0",x"80",x"00",x"00",x"3C",x"28",
    x"10",x"08",x"88",x"BF",x"00",x"3C",x"10",x"08",
    x"00",x"A0",x"80",x"02",x"00",x"00",x"C3",x"00",
    x"E3",x"3C",x"3C",x"10",x"10",x"10",x"10",x"36",
    x"08",x"08",x"8B",x"BF",x"00",x"29",x"00",x"A0",
    x"BF",x"2E",x"C7",x"E8",x"0C",x"20",x"3E",x"10",
    x"32",x"20",x"10",x"32",x"20",x"10",x"32",x"20",
    x"32",x"02",x"11",x"20",x"88",x"BF",x"0C",x"20",
    x"10",x"32",x"20",x"10",x"32",x"20",x"32",x"20",
    x"C3",x"00",x"E3",x"3E",x"10",x"36",x"0C",x"20",
    x"10",x"36",x"20",x"10",x"36",x"20",x"10",x"36",
    x"20",x"36",x"20",x"36",x"20",x"36",x"C7",x"E8",
    x"E3",x"3E",x"10",x"36",x"0C",x"20",x"10",x"36",
    x"20",x"10",x"36",x"20",x"10",x"36",x"20",x"16",
    x"3C",x"06",x"10",x"10",x"10",x"11",x"20",x"08",
    x"8A",x"BF",x"00",x"2B",x"8A",x"BF",x"00",x"11",
    x"88",x"BF",x"0C",x"20",x"10",x"36",x"20",x"10",
    x"36",x"20",x"36",x"20",x"C7",x"E8",x"E3",x"3C",
    x"10",x"10",x"28",x"10",x"28",x"10",x"28",x"10",
    x"28",x"10",x"28",x"28",x"28",x"10",x"28",x"28",
    x"10",x"28",x"10",x"28",x"10",x"10",x"10",x"28",
    x"3C",x"80",x"10",x"09",x"8B",x"BF",x"00",x"28",
    x"00",x"48",x"A0",x"BF",x"08",x"0C",x"10",x"0C",
    x"20",x"00",x"A0",x"BF",x"00",x"3C",x"3C",x"10",
    x"10",x"80",x"10",x"08",x"8B",x"BF",x"00",x"28",
    x"00",x"48",x"A1",x"BF",x"08",x"3C",x"3C",x"3C",
    x"3C",x"3C",x"3C",x"3C",x"3C",x"16",x"16",x"17",
    x"17",x"15",x"15",x"15",x"10",x"14",x"14",x"0C",
    x"88",x"BF",x"00",x"0D",x"08",x"A0",x"80",x"A0",
    x"3C",x"3C",x"10",x"10",x"80",x"10",x"08",x"8B",
    x"BF",x"00",x"28",x"00",x"48",x"A1",x"BF",x"08",
    x"C7",x"E8",x"80",x"A0",x"10",x"3E",x"00",x"00",
    x"A1",x"80",x"00",x"10",x"14",x"30",x"0D",x"0C",
    x"8B",x"BF",x"00",x"28",x"00",x"A0",x"BF",x"28",
    x"10",x"80",x"14",x"0C",x"89",x"BF",x"00",x"28",
    x"00",x"48",x"A0",x"BF",x"08",x"3C",x"14",x"80",
    x"10",x"A0",x"BF",x"00",x"3C",x"14",x"80",x"10",
    x"0C",x"89",x"BF",x"00",x"28",x"00",x"48",x"A0",
    x"BF",x"08",x"10",x"80",x"14",x"0C",x"89",x"BF",
    x"00",x"28",x"00",x"48",x"A0",x"BF",x"08",x"10",
    x"00",x"00",x"FF",x"10",x"FF",x"10",x"04",x"A4",
    x"BF",x"10",x"80",x"14",x"0C",x"89",x"BF",x"00",
    x"28",x"00",x"48",x"A0",x"BF",x"08",x"10",x"00",
    x"00",x"FF",x"10",x"04",x"A4",x"BF",x"00",x"10",
    x"04",x"80",x"0C",x"14",x"10",x"2A",x"04",x"FF",
    x"32",x"A4",x"BF",x"10",x"80",x"14",x"0C",x"89",
    x"BF",x"00",x"28",x"00",x"48",x"A0",x"BF",x"08",
    x"10",x"0C",x"3E",x"00",x"10",x"10",x"2B",x"2B",
    x"A3",x"80",x"00",x"10",x"14",x"30",x"0D",x"0C",
    x"8B",x"BF",x"00",x"28",x"00",x"A0",x"BF",x"28",
    x"10",x"80",x"14",x"0C",x"89",x"BF",x"00",x"28",
    x"00",x"48",x"A0",x"BF",x"08",x"3C",x"14",x"80",
    x"10",x"A0",x"BF",x"00",x"10",x"80",x"14",x"0C",
    x"89",x"BF",x"00",x"28",x"00",x"48",x"A0",x"BF",
    x"08",x"BF",x"0C",x"89",x"BF",x"00",x"28",x"00",
    x"48",x"A0",x"BF",x"08",x"BF",x"14",x"80",x"10",
    x"80",x"0C",x"89",x"BF",x"00",x"28",x"00",x"48",
    x"A0",x"BF",x"08",x"BF",x"0C",x"88",x"BF",x"3C",
    x"10",x"08",x"00",x"08",x"A0",x"BF",x"28",x"06",
    x"C0",x"00",x"0C",x"88",x"BF",x"00",x"0D",x"A0",
    x"BF",x"A0",x"BF",x"00",x"BF",x"0C",x"88",x"BF",
    x"00",x"0D",x"A0",x"BF",x"A0",x"BF",x"00",x"BF",
    x"FF",x"0C",x"FF",x"0A",x"06",x"27",x"10",x"FF",
    x"0A",x"2E",x"0A",x"06",x"80",x"06",x"FF",x"06",
    x"2C",x"04",x"07",x"A6",x"BF",x"00",x"80",x"00",
    x"FF",x"00",x"FF",x"0A",x"0A",x"FF",x"2A",x"06",
    x"0A",x"FF",x"27",x"04",x"0A",x"2E",x"3F",x"06",
    x"0C",x"2E",x"10",x"80",x"06",x"FF",x"06",x"2C",
    x"04",x"07",x"A6",x"BF",x"00",x"80",x"00",x"FF",
    x"00",x"FF",x"0A",x"FF",x"0A",x"0A",x"2C",x"FF",
    x"04",x"2C",x"06",x"0A",x"FF",x"27",x"04",x"0A",
    x"2E",x"3F",x"06",x"0C",x"2E",x"10",x"80",x"06",
    x"FF",x"06",x"2C",x"04",x"07",x"A6",x"BF",x"00",
    x"00",x"A4",x"80",x"10",x"FF",x"00",x"BF",x"00",
    x"6F",x"6F",x"72",x"00",x"0A",x"00",x"58",x"52",
    x"0D",x"00",x"0D",x"00",x"4F",x"4C",x"20",x"52",
    x"0A",x"00",x"4C",x"0A",x"4C",x"20",x"54",x"00",
    x"4C",x"20",x"54",x"00",x"45",x"45",x"52",x"00",
    x"45",x"4F",x"00",x"00",x"00",x"00",x"31",x"35",
    x"39",x"44",x"10",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );

  CONSTANT INIT5_2 : type_mem:=(
    x"00",x"62",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"00",x"E2",x"00",x"00",
    x"00",x"E3",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"00",x"00",x"40",x"80",x"00",x"00",x"40",x"80",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"00",x"60",x"60",x"20",x"00",x"40",x"C0",x"21",
    x"80",x"20",x"22",x"80",x"20",x"20",x"80",x"00",
    x"00",x"00",x"00",x"63",x"00",x"00",x"20",x"80",
    x"80",x"00",x"A3",x"00",x"E3",x"00",x"00",x"01",
    x"00",x"00",x"00",x"20",x"40",x"24",x"00",x"00",
    x"00",x"00",x"00",x"00",x"40",x"00",x"40",x"00",
    x"00",x"20",x"20",x"00",x"00",x"40",x"00",x"00",
    x"00",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",
    x"A0",x"00",x"00",x"40",x"80",x"00",x"00",x"00",
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",
    x"A0",x"00",x"00",x"40",x"80",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"0C",x"0D",x"0D",x"0E",x"08",x"08",x"08",x"0D",
    x"00",x"E0",x"00",x"00",x"E0",x"00",x"00",x"E0",
    x"00",x"00",x"E0",x"00",x"00",x"E0",x"00",x"00",
    x"E0",x"00",x"44",x"60",x"40",x"A0",x"FF",x"00",
    x"44",x"60",x"40",x"E0",x"00",x"44",x"60",x"00",
    x"60",x"40",x"20",x"FF",x"00",x"80",x"20",x"00",
    x"E0",x"FF",x"00",x"E0",x"00",x"44",x"60",x"40",
    x"A0",x"FF",x"00",x"44",x"60",x"40",x"E0",x"00",
    x"20",x"44",x"60",x"40",x"20",x"40",x"20",x"40",
    x"20",x"40",x"20",x"40",x"40",x"40",x"20",x"40",
    x"40",x"3F",x"40",x"20",x"40",x"3F",x"40",x"E0",
    x"00",x"44",x"60",x"40",x"A0",x"FF",x"00",x"44",
    x"60",x"40",x"60",x"00",x"7F",x"7F",x"44",x"A0",
    x"60",x"40",x"E0",x"FF",x"00",x"44",x"60",x"40",
    x"7F",x"60",x"00",x"00",x"7F",x"40",x"E0",x"00",
    x"BF",x"44",x"00",x"A0",x"E3",x"20",x"A0",x"20",
    x"C0",x"80",x"20",x"FF",x"00",x"00",x"60",x"60",
    x"FF",x"20",x"E0",x"00",x"3C",x"40",x"40",x"20",
    x"00",x"40",x"20",x"00",x"40",x"20",x"00",x"40",
    x"00",x"00",x"00",x"40",x"E0",x"FF",x"3C",x"C0",
    x"20",x"00",x"C0",x"20",x"00",x"C0",x"00",x"C0",
    x"E0",x"00",x"BF",x"40",x"20",x"00",x"3C",x"80",
    x"20",x"00",x"80",x"20",x"00",x"80",x"20",x"00",
    x"80",x"00",x"80",x"00",x"80",x"00",x"E0",x"00",
    x"BF",x"40",x"20",x"00",x"3C",x"80",x"20",x"00",
    x"80",x"20",x"00",x"80",x"20",x"00",x"80",x"00",
    x"44",x"00",x"E0",x"20",x"E0",x"00",x"80",x"C0",
    x"A0",x"FF",x"00",x"00",x"E0",x"FF",x"00",x"00",
    x"A0",x"FF",x"3C",x"80",x"20",x"00",x"80",x"20",
    x"00",x"80",x"00",x"80",x"E0",x"00",x"BF",x"44",
    x"20",x"A0",x"40",x"20",x"40",x"20",x"40",x"20",
    x"40",x"20",x"40",x"40",x"40",x"20",x"40",x"40",
    x"3F",x"40",x"20",x"40",x"00",x"3F",x"A0",x"40",
    x"00",x"00",x"62",x"00",x"60",x"FF",x"00",x"80",
    x"60",x"40",x"E0",x"FF",x"40",x"00",x"3F",x"04",
    x"40",x"60",x"40",x"FF",x"00",x"44",x"00",x"A0",
    x"62",x"00",x"A0",x"80",x"60",x"FF",x"00",x"C0",
    x"60",x"40",x"20",x"FF",x"40",x"44",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"A0",x"E3",x"23",
    x"63",x"E3",x"A3",x"62",x"20",x"60",x"60",x"00",
    x"60",x"FF",x"00",x"00",x"60",x"60",x"00",x"60",
    x"44",x"00",x"A0",x"62",x"00",x"A0",x"80",x"60",
    x"FF",x"00",x"C0",x"60",x"40",x"20",x"FF",x"40",
    x"E0",x"00",x"00",x"60",x"20",x"40",x"04",x"40",
    x"3F",x"00",x"60",x"20",x"60",x"60",x"80",x"00",
    x"60",x"FF",x"00",x"C0",x"A0",x"A0",x"FF",x"60",
    x"00",x"00",x"60",x"00",x"20",x"FF",x"00",x"80",
    x"60",x"40",x"E0",x"FF",x"40",x"00",x"60",x"00",
    x"62",x"40",x"FF",x"00",x"00",x"60",x"00",x"63",
    x"00",x"20",x"FF",x"00",x"80",x"60",x"40",x"E0",
    x"FF",x"40",x"00",x"00",x"60",x"00",x"20",x"FF",
    x"00",x"80",x"60",x"40",x"E0",x"FF",x"40",x"20",
    x"00",x"04",x"FF",x"00",x"FF",x"00",x"C0",x"C0",
    x"FF",x"00",x"00",x"60",x"00",x"20",x"FF",x"00",
    x"80",x"60",x"40",x"E0",x"FF",x"40",x"20",x"00",
    x"04",x"FE",x"00",x"C0",x"C0",x"FF",x"00",x"20",
    x"A0",x"00",x"00",x"C0",x"00",x"60",x"E0",x"FE",
    x"60",x"C0",x"FF",x"00",x"00",x"60",x"00",x"20",
    x"FF",x"00",x"80",x"60",x"40",x"E0",x"FF",x"40",
    x"20",x"00",x"40",x"04",x"40",x"40",x"60",x"20",
    x"00",x"00",x"60",x"20",x"60",x"60",x"80",x"00",
    x"60",x"FF",x"00",x"C0",x"A0",x"A0",x"FF",x"60",
    x"00",x"00",x"60",x"00",x"20",x"FF",x"00",x"80",
    x"60",x"40",x"E0",x"FF",x"40",x"00",x"60",x"00",
    x"63",x"40",x"FF",x"00",x"00",x"00",x"60",x"00",
    x"20",x"FF",x"00",x"80",x"60",x"40",x"E0",x"FF",
    x"40",x"FF",x"00",x"20",x"FF",x"00",x"80",x"60",
    x"40",x"E0",x"FF",x"40",x"FF",x"60",x"00",x"00",
    x"00",x"00",x"20",x"FF",x"00",x"80",x"60",x"40",
    x"E0",x"FF",x"40",x"FF",x"00",x"60",x"FF",x"44",
    x"60",x"40",x"7F",x"60",x"60",x"FF",x"60",x"80",
    x"40",x"00",x"00",x"60",x"FF",x"00",x"00",x"60",
    x"FE",x"60",x"FF",x"00",x"FE",x"00",x"60",x"FF",
    x"00",x"00",x"60",x"FE",x"60",x"FF",x"00",x"FE",
    x"FE",x"00",x"FE",x"20",x"3F",x"BF",x"20",x"FE",
    x"20",x"20",x"20",x"00",x"00",x"00",x"FD",x"60",
    x"C0",x"E0",x"BF",x"40",x"FF",x"00",x"00",x"40",
    x"FD",x"00",x"FD",x"20",x"20",x"FD",x"20",x"7F",
    x"20",x"FD",x"BF",x"C0",x"20",x"20",x"C0",x"00",
    x"00",x"00",x"20",x"00",x"00",x"FD",x"60",x"C0",
    x"E0",x"BF",x"40",x"FF",x"00",x"00",x"40",x"FD",
    x"00",x"FD",x"20",x"FD",x"20",x"20",x"E0",x"FD",
    x"C0",x"E0",x"7F",x"20",x"FD",x"BF",x"C0",x"20",
    x"20",x"C0",x"00",x"00",x"00",x"20",x"00",x"00",
    x"FD",x"60",x"C0",x"E0",x"BF",x"40",x"FF",x"00",
    x"40",x"80",x"00",x"00",x"FD",x"00",x"FE",x"00",
    x"6F",x"61",x"0A",x"00",x"0D",x"00",x"45",x"41",
    x"00",x"00",x"00",x"00",x"54",x"41",x"3A",x"41",
    x"0D",x"00",x"41",x"0D",x"41",x"57",x"45",x"00",
    x"41",x"54",x"0A",x"00",x"53",x"52",x"0A",x"00",
    x"53",x"4B",x"00",x"00",x"00",x"00",x"32",x"36",
    x"41",x"45",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );

  CONSTANT INIT5_3 : type_mem:=(
    x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",
    x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",
    x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"04",x"A0",x"00",x"02",x"00",x"00",x"00",x"00",
    x"80",x"03",x"00",x"80",x"01",x"00",x"80",x"00",
    x"00",x"00",x"04",x"00",x"01",x"0E",x"00",x"00",
    x"00",x"03",x"78",x"03",x"78",x"00",x"00",x"4F",
    x"00",x"00",x"00",x"9E",x"00",x"00",x"60",x"00",
    x"00",x"00",x"00",x"08",x"00",x"08",x"00",x"00",
    x"01",x"01",x"07",x"01",x"00",x"00",x"00",x"00",
    x"00",x"00",x"08",x"10",x"18",x"20",x"28",x"30",
    x"38",x"00",x"13",x"00",x"00",x"00",x"00",x"00",
    x"01",x"07",x"13",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"08",x"10",x"18",x"20",x"28",x"30",
    x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"1E",x"1E",x"1E",x"1E",
    x"9E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",
    x"E8",x"40",x"A0",x"1C",x"FC",x"FC",x"FC",x"14",
    x"00",x"08",x"00",x"00",x"08",x"00",x"00",x"08",
    x"00",x"00",x"08",x"00",x"00",x"08",x"00",x"00",
    x"08",x"00",x"00",x"04",x"00",x"04",x"FE",x"00",
    x"00",x"06",x"00",x"08",x"00",x"00",x"06",x"08",
    x"04",x"00",x"04",x"FE",x"00",x"00",x"01",x"00",
    x"00",x"F8",x"00",x"08",x"00",x"00",x"04",x"00",
    x"01",x"FE",x"00",x"00",x"06",x"00",x"08",x"00",
    x"04",x"00",x"04",x"00",x"44",x"00",x"0C",x"00",
    x"0E",x"00",x"0D",x"00",x"00",x"00",x"03",x"00",
    x"00",x"C1",x"00",x"05",x"00",x"EA",x"00",x"08",
    x"00",x"00",x"04",x"00",x"01",x"FE",x"00",x"00",
    x"06",x"00",x"40",x"03",x"D0",x"C9",x"00",x"04",
    x"04",x"00",x"01",x"FE",x"00",x"00",x"06",x"00",
    x"C9",x"40",x"04",x"02",x"D0",x"02",x"08",x"00",
    x"A0",x"00",x"03",x"06",x"58",x"00",x"04",x"1C",
    x"0D",x"00",x"04",x"FE",x"00",x"00",x"01",x"08",
    x"F7",x"04",x"08",x"00",x"00",x"00",x"00",x"50",
    x"02",x"00",x"FF",x"02",x"00",x"40",x"02",x"00",
    x"02",x"02",x"00",x"00",x"80",x"FD",x"00",x"00",
    x"FF",x"02",x"00",x"50",x"02",x"00",x"02",x"00",
    x"08",x"00",x"A0",x"00",x"50",x"01",x"00",x"00",
    x"FF",x"01",x"00",x"60",x"01",x"00",x"D0",x"01",
    x"00",x"01",x"00",x"01",x"00",x"01",x"08",x"00",
    x"A0",x"00",x"50",x"01",x"00",x"00",x"FF",x"01",
    x"00",x"20",x"01",x"00",x"D0",x"01",x"00",x"01",
    x"00",x"01",x"06",x"2D",x"04",x"00",x"00",x"00",
    x"04",x"FE",x"00",x"00",x"80",x"F8",x"00",x"00",
    x"80",x"FE",x"00",x"00",x"FF",x"01",x"00",x"50",
    x"01",x"00",x"01",x"00",x"08",x"00",x"98",x"00",
    x"04",x"04",x"00",x"44",x"00",x"0C",x"00",x"0E",
    x"00",x"0D",x"00",x"00",x"00",x"03",x"00",x"00",
    x"C1",x"00",x"05",x"00",x"01",x"EA",x"06",x"00",
    x"03",x"08",x"C0",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"00",x"FF",x"00",
    x"00",x"04",x"02",x"FD",x"00",x"00",x"03",x"06",
    x"D0",x"08",x"04",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"00",x"01",x"03",
    x"03",x"03",x"03",x"03",x"03",x"00",x"50",x"10",
    x"20",x"40",x"58",x"E8",x"00",x"04",x"06",x"00",
    x"01",x"FE",x"00",x"00",x"5F",x"58",x"14",x"57",
    x"00",x"03",x"06",x"D8",x"08",x"04",x"00",x"04",
    x"FE",x"00",x"00",x"01",x"00",x"00",x"F8",x"00",
    x"08",x"00",x"C3",x"53",x"00",x"00",x"00",x"03",
    x"FF",x"20",x"04",x"00",x"06",x"1C",x"04",x"00",
    x"04",x"FE",x"00",x"00",x"01",x"08",x"F7",x"04",
    x"15",x"08",x"06",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"03",x"06",x"1C",
    x"F0",x"02",x"DD",x"00",x"03",x"06",x"08",x"08",
    x"00",x"04",x"FE",x"00",x"00",x"01",x"00",x"00",
    x"F8",x"00",x"1C",x"1F",x"06",x"00",x"04",x"FE",
    x"00",x"00",x"01",x"00",x"00",x"F8",x"00",x"00",
    x"80",x"00",x"08",x"13",x"1C",x"13",x"18",x"19",
    x"FA",x"1C",x"08",x"06",x"00",x"04",x"FE",x"00",
    x"00",x"01",x"00",x"00",x"F8",x"00",x"00",x"80",
    x"00",x"F1",x"13",x"18",x"19",x"FC",x"00",x"00",
    x"02",x"08",x"00",x"19",x"13",x"10",x"02",x"C5",
    x"10",x"18",x"F9",x"1D",x"08",x"06",x"00",x"04",
    x"FE",x"00",x"00",x"01",x"00",x"00",x"F8",x"00",
    x"00",x"00",x"00",x"00",x"04",x"03",x"10",x"10",
    x"0D",x"20",x"02",x"00",x"06",x"1C",x"04",x"00",
    x"04",x"FE",x"00",x"00",x"01",x"08",x"F7",x"04",
    x"15",x"08",x"06",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"03",x"06",x"19",
    x"30",x"02",x"DA",x"00",x"17",x"08",x"06",x"00",
    x"04",x"FE",x"00",x"00",x"01",x"00",x"00",x"F8",
    x"00",x"2E",x"00",x"04",x"FE",x"00",x"00",x"01",
    x"00",x"00",x"F8",x"00",x"23",x"06",x"09",x"1B",
    x"0C",x"00",x"04",x"FE",x"00",x"00",x"01",x"00",
    x"00",x"F8",x"00",x"14",x"00",x"01",x"FE",x"00",
    x"06",x"00",x"D0",x"FF",x"07",x"0A",x"02",x"01",
    x"00",x"00",x"00",x"01",x"FE",x"00",x"00",x"0D",
    x"FF",x"0A",x"F8",x"00",x"FB",x"00",x"01",x"FE",
    x"00",x"00",x"0D",x"F4",x"0A",x"F8",x"00",x"F0",
    x"09",x"00",x"07",x"FF",x"FD",x"FC",x"00",x"02",
    x"FF",x"08",x"FF",x"08",x"06",x"13",x"FB",x"01",
    x"00",x"01",x"FC",x"01",x"FA",x"00",x"43",x"18",
    x"F1",x"00",x"EF",x"FF",x"FF",x"EC",x"08",x"FC",
    x"FF",x"E8",x"FC",x"18",x"FF",x"08",x"00",x"08",
    x"00",x"01",x"00",x"06",x"13",x"DC",x"01",x"00",
    x"01",x"FC",x"01",x"FA",x"00",x"24",x"18",x"D2",
    x"00",x"D0",x"FF",x"CE",x"FF",x"FF",x"08",x"CA",
    x"08",x"08",x"FB",x"FF",x"C5",x"FC",x"18",x"FF",
    x"08",x"00",x"08",x"00",x"01",x"00",x"06",x"13",
    x"B9",x"01",x"00",x"01",x"FC",x"01",x"FA",x"00",
    x"18",x"18",x"02",x"18",x"AD",x"00",x"91",x"00",
    x"74",x"64",x"0D",x"00",x"00",x"00",x"43",x"4D",
    x"00",x"00",x"00",x"00",x"20",x"4E",x"20",x"53",
    x"00",x"00",x"4E",x"00",x"53",x"52",x"0A",x"00",
    x"53",x"45",x"0D",x"00",x"54",x"52",x"0D",x"00",
    x"54",x"0A",x"00",x"00",x"00",x"00",x"33",x"37",
    x"42",x"46",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );


  CONSTANT INIT20_0 : type_mem:=(
    x"03",x"81",x"01",x"FF",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"27",x"81",x"A1",x"01",
    x"27",x"81",x"A1",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"01",x"01",x"81",x"81",x"01",x"01",x"81",x"81",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"03",x"82",x"81",x"81",x"03",x"81",x"03",x"84",
    x"C2",x"82",x"84",x"C2",x"82",x"84",x"C2",x"01",
    x"01",x"01",x"03",x"82",x"9C",x"BC",x"A0",x"E0",
    x"C1",x"05",x"84",x"07",x"86",x"82",x"01",x"40",
    x"01",x"01",x"03",x"84",x"C4",x"82",x"C2",x"01",
    x"01",x"81",x"01",x"03",x"81",x"03",x"81",x"01",
    x"A6",x"83",x"A1",x"82",x"81",x"81",x"01",x"01",
    x"01",x"E0",x"E4",x"E8",x"EC",x"F0",x"F4",x"F8",
    x"FC",x"81",x"82",x"81",x"81",x"01",x"01",x"01",
    x"A7",x"A1",x"A0",x"81",x"01",x"01",x"01",x"81",
    x"81",x"E0",x"E4",x"E8",x"EC",x"F0",x"F4",x"F8",
    x"FC",x"81",x"81",x"81",x"81",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"91",x"01",x"01",x"01",
    x"91",x"01",x"01",x"01",x"F0",x"FD",x"FE",x"EF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"D0",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
    x"D2",x"81",x"01",x"D2",x"81",x"01",x"D2",x"81",
    x"01",x"D0",x"81",x"01",x"D0",x"81",x"01",x"D0",
    x"81",x"01",x"03",x"82",x"C4",x"80",x"02",x"01",
    x"03",x"82",x"D0",x"81",x"01",x"03",x"84",x"10",
    x"82",x"C8",x"80",x"02",x"01",x"C6",x"90",x"C6",
    x"80",x"12",x"C6",x"81",x"01",x"03",x"82",x"C4",
    x"80",x"02",x"01",x"03",x"82",x"D0",x"81",x"01",
    x"84",x"03",x"82",x"C4",x"84",x"C4",x"84",x"C4",
    x"84",x"C4",x"86",x"C6",x"C0",x"C4",x"84",x"C4",
    x"C4",x"84",x"C4",x"84",x"C4",x"84",x"C4",x"81",
    x"01",x"03",x"82",x"C4",x"80",x"02",x"01",x"03",
    x"82",x"C2",x"80",x"08",x"84",x"84",x"03",x"85",
    x"82",x"C6",x"80",x"02",x"01",x"03",x"82",x"C2",
    x"90",x"80",x"18",x"90",x"82",x"90",x"81",x"01",
    x"9D",x"05",x"07",x"88",x"86",x"82",x"84",x"9B",
    x"DA",x"D8",x"80",x"02",x"01",x"DA",x"82",x"80",
    x"12",x"B1",x"81",x"81",x"03",x"C0",x"05",x"86",
    x"C6",x"C0",x"86",x"C6",x"C0",x"86",x"C6",x"C0",
    x"D2",x"88",x"C6",x"C0",x"80",x"02",x"07",x"C0",
    x"82",x"C2",x"C0",x"88",x"C8",x"C0",x"C2",x"C0",
    x"81",x"01",x"9D",x"03",x"88",x"C8",x"05",x"C0",
    x"86",x"C6",x"C0",x"9A",x"DA",x"C0",x"9A",x"DA",
    x"C0",x"C6",x"C0",x"C8",x"C0",x"C6",x"81",x"81",
    x"9D",x"03",x"84",x"C4",x"05",x"C0",x"86",x"C6",
    x"C0",x"86",x"C6",x"C0",x"86",x"C6",x"C0",x"C6",
    x"07",x"88",x"98",x"9A",x"86",x"D6",x"C0",x"D4",
    x"80",x"02",x"01",x"DA",x"80",x"02",x"01",x"C4",
    x"80",x"02",x"05",x"C0",x"86",x"C6",x"C0",x"88",
    x"C8",x"C0",x"C6",x"C0",x"81",x"81",x"9D",x"05",
    x"86",x"82",x"C6",x"86",x"C6",x"86",x"C6",x"86",
    x"C6",x"88",x"C8",x"C0",x"C6",x"86",x"C6",x"C6",
    x"86",x"C6",x"86",x"C6",x"88",x"86",x"84",x"C6",
    x"03",x"10",x"82",x"DA",x"80",x"02",x"01",x"C6",
    x"82",x"C6",x"80",x"12",x"C6",x"03",x"86",x"05",
    x"C6",x"82",x"80",x"12",x"01",x"05",x"03",x"86",
    x"82",x"10",x"84",x"DA",x"80",x"02",x"01",x"C8",
    x"82",x"C8",x"80",x"12",x"C8",x"23",x"35",x"37",
    x"39",x"3B",x"2F",x"2D",x"2B",x"B4",x"B6",x"B8",
    x"BA",x"AE",x"AC",x"AA",x"A4",x"A0",x"A8",x"C2",
    x"80",x"02",x"01",x"C2",x"82",x"80",x"12",x"80",
    x"05",x"03",x"86",x"82",x"10",x"84",x"DA",x"80",
    x"02",x"01",x"C8",x"82",x"C8",x"80",x"12",x"C8",
    x"81",x"81",x"12",x"80",x"82",x"07",x"05",x"C8",
    x"80",x"22",x"82",x"84",x"86",x"89",x"C8",x"DA",
    x"80",x"02",x"01",x"C8",x"84",x"80",x"32",x"83",
    x"82",x"10",x"84",x"C8",x"80",x"02",x"01",x"C6",
    x"82",x"C6",x"80",x"12",x"C6",x"03",x"84",x"10",
    x"82",x"80",x"12",x"01",x"03",x"84",x"10",x"82",
    x"C8",x"80",x"02",x"01",x"C6",x"82",x"C6",x"80",
    x"12",x"C6",x"82",x"10",x"84",x"C8",x"80",x"02",
    x"01",x"C6",x"82",x"C6",x"80",x"12",x"C6",x"A6",
    x"31",x"33",x"7F",x"90",x"7F",x"90",x"A6",x"80",
    x"12",x"82",x"10",x"84",x"C8",x"80",x"02",x"01",
    x"C6",x"82",x"C6",x"80",x"12",x"C6",x"A6",x"31",
    x"33",x"7F",x"90",x"A6",x"80",x"12",x"01",x"A6",
    x"B0",x"10",x"33",x"D2",x"90",x"93",x"A6",x"7F",
    x"93",x"80",x"0A",x"82",x"10",x"84",x"C8",x"80",
    x"02",x"01",x"C6",x"82",x"C6",x"80",x"12",x"C6",
    x"82",x"09",x"07",x"05",x"DA",x"D8",x"9B",x"99",
    x"80",x"22",x"82",x"84",x"86",x"89",x"C8",x"DA",
    x"80",x"02",x"01",x"C8",x"84",x"80",x"32",x"83",
    x"82",x"10",x"84",x"C8",x"80",x"02",x"01",x"C6",
    x"82",x"C6",x"80",x"12",x"C6",x"03",x"84",x"10",
    x"82",x"80",x"12",x"01",x"82",x"10",x"84",x"C8",
    x"80",x"02",x"01",x"C6",x"82",x"C6",x"80",x"12",
    x"C6",x"30",x"C8",x"80",x"02",x"01",x"C6",x"82",
    x"C6",x"80",x"12",x"C6",x"30",x"84",x"12",x"82",
    x"30",x"C8",x"80",x"02",x"01",x"C6",x"82",x"C6",
    x"80",x"12",x"C6",x"30",x"C2",x"80",x"02",x"03",
    x"82",x"C2",x"82",x"82",x"80",x"18",x"83",x"C2",
    x"81",x"01",x"C2",x"80",x"02",x"01",x"C2",x"80",
    x"02",x"80",x"12",x"01",x"30",x"C2",x"80",x"02",
    x"01",x"C2",x"80",x"02",x"80",x"12",x"01",x"30",
    x"7F",x"27",x"7F",x"B0",x"B0",x"F0",x"B2",x"7F",
    x"B0",x"B1",x"90",x"B0",x"10",x"A6",x"7F",x"B2",
    x"D0",x"A6",x"C2",x"80",x"0A",x"01",x"10",x"B0",
    x"7F",x"01",x"7F",x"B2",x"90",x"7F",x"A7",x"B2",
    x"B0",x"7F",x"F2",x"B0",x"90",x"B1",x"03",x"B0",
    x"27",x"B0",x"B2",x"10",x"A6",x"7F",x"B2",x"D0",
    x"A6",x"C2",x"80",x"0A",x"01",x"10",x"B0",x"7F",
    x"01",x"7F",x"B2",x"7F",x"A6",x"90",x"A7",x"7F",
    x"A6",x"A7",x"B2",x"B0",x"7F",x"F2",x"B0",x"90",
    x"B1",x"03",x"B0",x"27",x"B0",x"B2",x"10",x"A6",
    x"7F",x"B2",x"D0",x"A6",x"C2",x"80",x"0A",x"01",
    x"B0",x"80",x"2A",x"A4",x"7F",x"01",x"30",x"00",
    x"42",x"6C",x"65",x"00",x"3E",x"00",x"45",x"20",
    x"0A",x"00",x"0A",x"00",x"4E",x"42",x"4B",x"45",
    x"45",x"00",x"42",x"4B",x"46",x"48",x"49",x"0D",
    x"46",x"48",x"53",x"00",x"54",x"20",x"4F",x"00",
    x"54",x"20",x"0D",x"00",x"3E",x"00",x"30",x"34",
    x"38",x"43",x"00",x"30",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );

  CONSTANT INIT20_1 : type_mem:=(
    x"3C",x"C0",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"3C",x"C4",x"50",x"00",
    x"3C",x"C4",x"50",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"00",x"10",x"20",x"30",x"40",x"50",x"60",x"70",
    x"80",x"90",x"A0",x"B0",x"C0",x"D0",x"E0",x"F0",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"00",x"00",x"C4",x"CC",x"00",x"00",x"C4",x"CC",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"00",x"10",x"88",x"90",x"3C",x"98",x"3F",x"10",
    x"A0",x"10",x"10",x"A0",x"10",x"10",x"A0",x"00",
    x"00",x"00",x"3C",x"10",x"10",x"10",x"10",x"23",
    x"0B",x"3C",x"10",x"3C",x"10",x"10",x"00",x"00",
    x"00",x"00",x"3C",x"10",x"20",x"10",x"A0",x"00",
    x"00",x"C0",x"00",x"3C",x"98",x"00",x"C0",x"00",
    x"10",x"34",x"2C",x"14",x"E0",x"90",x"00",x"00",
    x"00",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",x"3B",
    x"3B",x"E8",x"10",x"C4",x"CC",x"00",x"00",x"00",
    x"2C",x"34",x"14",x"94",x"00",x"00",x"00",x"E8",
    x"E8",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",
    x"1B",x"E0",x"E0",x"C4",x"CC",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"D0",x"00",x"00",x"00",
    x"D0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"10",x"20",x"30",x"40",x"50",x"60",x"70",
    x"00",x"00",x"A0",x"B0",x"C0",x"D0",x"E0",x"F0",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"2A",x"C3",x"00",x"32",x"C3",x"00",x"22",x"C3",
    x"00",x"0A",x"C3",x"00",x"12",x"C3",x"00",x"02",
    x"C3",x"00",x"3C",x"10",x"08",x"88",x"BF",x"00",
    x"3C",x"10",x"28",x"C3",x"00",x"3C",x"10",x"80",
    x"10",x"08",x"89",x"BF",x"00",x"28",x"02",x"4A",
    x"A0",x"BF",x"0A",x"C3",x"00",x"3C",x"10",x"08",
    x"88",x"BF",x"00",x"3C",x"10",x"08",x"C3",x"00",
    x"10",x"3C",x"10",x"28",x"10",x"28",x"10",x"28",
    x"10",x"28",x"10",x"28",x"28",x"28",x"10",x"28",
    x"28",x"10",x"28",x"10",x"28",x"10",x"28",x"C3",
    x"00",x"3C",x"10",x"08",x"88",x"BF",x"00",x"3C",
    x"10",x"08",x"A0",x"80",x"00",x"00",x"3C",x"28",
    x"10",x"08",x"88",x"BF",x"00",x"3C",x"10",x"08",
    x"00",x"A0",x"80",x"02",x"00",x"00",x"C3",x"00",
    x"E3",x"3C",x"3C",x"10",x"10",x"10",x"10",x"36",
    x"08",x"08",x"8B",x"BF",x"00",x"29",x"00",x"A0",
    x"BF",x"2E",x"C7",x"E8",x"0C",x"20",x"3E",x"10",
    x"32",x"20",x"10",x"32",x"20",x"10",x"32",x"20",
    x"32",x"02",x"11",x"20",x"88",x"BF",x"0C",x"20",
    x"10",x"32",x"20",x"10",x"32",x"20",x"32",x"20",
    x"C3",x"00",x"E3",x"3E",x"10",x"36",x"0C",x"20",
    x"10",x"36",x"20",x"10",x"36",x"20",x"10",x"36",
    x"20",x"36",x"20",x"36",x"20",x"36",x"C7",x"E8",
    x"E3",x"3E",x"10",x"36",x"0C",x"20",x"10",x"36",
    x"20",x"10",x"36",x"20",x"10",x"36",x"20",x"16",
    x"3C",x"06",x"10",x"10",x"10",x"11",x"20",x"08",
    x"8A",x"BF",x"00",x"2B",x"8A",x"BF",x"00",x"11",
    x"88",x"BF",x"0C",x"20",x"10",x"36",x"20",x"10",
    x"36",x"20",x"36",x"20",x"C7",x"E8",x"E3",x"3C",
    x"10",x"10",x"28",x"10",x"28",x"10",x"28",x"10",
    x"28",x"10",x"28",x"28",x"28",x"10",x"28",x"28",
    x"10",x"28",x"10",x"28",x"10",x"10",x"10",x"28",
    x"3C",x"80",x"10",x"09",x"8B",x"BF",x"00",x"28",
    x"00",x"48",x"A0",x"BF",x"08",x"0C",x"10",x"0C",
    x"20",x"00",x"A0",x"BF",x"00",x"3C",x"3C",x"10",
    x"10",x"80",x"10",x"08",x"8B",x"BF",x"00",x"28",
    x"00",x"48",x"A1",x"BF",x"08",x"3C",x"3C",x"3C",
    x"3C",x"3C",x"3C",x"3C",x"3C",x"16",x"16",x"17",
    x"17",x"15",x"15",x"15",x"10",x"14",x"14",x"0C",
    x"88",x"BF",x"00",x"0D",x"08",x"A0",x"80",x"A0",
    x"3C",x"3C",x"10",x"10",x"80",x"10",x"08",x"8B",
    x"BF",x"00",x"28",x"00",x"48",x"A1",x"BF",x"08",
    x"C7",x"E8",x"80",x"A0",x"10",x"3E",x"00",x"00",
    x"A1",x"80",x"00",x"10",x"14",x"30",x"0D",x"0C",
    x"8B",x"BF",x"00",x"28",x"00",x"A0",x"BF",x"28",
    x"10",x"80",x"14",x"0C",x"89",x"BF",x"00",x"28",
    x"00",x"48",x"A0",x"BF",x"08",x"3C",x"14",x"80",
    x"10",x"A0",x"BF",x"00",x"3C",x"14",x"80",x"10",
    x"0C",x"89",x"BF",x"00",x"28",x"00",x"48",x"A0",
    x"BF",x"08",x"10",x"80",x"14",x"0C",x"89",x"BF",
    x"00",x"28",x"00",x"48",x"A0",x"BF",x"08",x"10",
    x"00",x"00",x"FF",x"10",x"FF",x"10",x"04",x"A4",
    x"BF",x"10",x"80",x"14",x"0C",x"89",x"BF",x"00",
    x"28",x"00",x"48",x"A0",x"BF",x"08",x"10",x"00",
    x"00",x"FF",x"10",x"04",x"A4",x"BF",x"00",x"10",
    x"04",x"80",x"0C",x"14",x"10",x"2A",x"04",x"FF",
    x"32",x"A4",x"BF",x"10",x"80",x"14",x"0C",x"89",
    x"BF",x"00",x"28",x"00",x"48",x"A0",x"BF",x"08",
    x"10",x"0C",x"3E",x"00",x"10",x"10",x"2B",x"2B",
    x"A3",x"80",x"00",x"10",x"14",x"30",x"0D",x"0C",
    x"8B",x"BF",x"00",x"28",x"00",x"A0",x"BF",x"28",
    x"10",x"80",x"14",x"0C",x"89",x"BF",x"00",x"28",
    x"00",x"48",x"A0",x"BF",x"08",x"3C",x"14",x"80",
    x"10",x"A0",x"BF",x"00",x"10",x"80",x"14",x"0C",
    x"89",x"BF",x"00",x"28",x"00",x"48",x"A0",x"BF",
    x"08",x"BF",x"0C",x"89",x"BF",x"00",x"28",x"00",
    x"48",x"A0",x"BF",x"08",x"BF",x"14",x"80",x"10",
    x"80",x"0C",x"89",x"BF",x"00",x"28",x"00",x"48",
    x"A0",x"BF",x"08",x"BF",x"0C",x"88",x"BF",x"3C",
    x"10",x"08",x"00",x"08",x"A0",x"BF",x"28",x"06",
    x"C0",x"00",x"0C",x"88",x"BF",x"00",x"0D",x"A0",
    x"BF",x"A0",x"BF",x"00",x"BF",x"0C",x"88",x"BF",
    x"00",x"0D",x"A0",x"BF",x"A0",x"BF",x"00",x"BF",
    x"FF",x"0C",x"FF",x"0A",x"06",x"27",x"10",x"FF",
    x"0A",x"2E",x"0A",x"06",x"80",x"06",x"FF",x"06",
    x"2C",x"04",x"07",x"A6",x"BF",x"00",x"80",x"00",
    x"FF",x"00",x"FF",x"0A",x"0A",x"FF",x"2A",x"06",
    x"0A",x"FF",x"27",x"04",x"0A",x"2E",x"3F",x"06",
    x"0C",x"2E",x"10",x"80",x"06",x"FF",x"06",x"2C",
    x"04",x"07",x"A6",x"BF",x"00",x"80",x"00",x"FF",
    x"00",x"FF",x"0A",x"FF",x"0A",x"0A",x"2C",x"FF",
    x"04",x"2C",x"06",x"0A",x"FF",x"27",x"04",x"0A",
    x"2E",x"3F",x"06",x"0C",x"2E",x"10",x"80",x"06",
    x"FF",x"06",x"2C",x"04",x"07",x"A6",x"BF",x"00",
    x"00",x"A4",x"80",x"10",x"FF",x"00",x"BF",x"00",
    x"6F",x"6F",x"72",x"00",x"0A",x"00",x"58",x"52",
    x"0D",x"00",x"0D",x"00",x"4F",x"4C",x"20",x"52",
    x"0A",x"00",x"4C",x"0A",x"4C",x"20",x"54",x"00",
    x"4C",x"20",x"54",x"00",x"45",x"45",x"52",x"00",
    x"45",x"4F",x"00",x"00",x"00",x"00",x"31",x"35",
    x"39",x"44",x"10",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );

  CONSTANT INIT20_2 : type_mem:=(
    x"00",x"62",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"00",x"E2",x"00",x"00",
    x"00",x"E3",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"00",x"00",x"40",x"80",x"00",x"00",x"40",x"80",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"00",x"60",x"60",x"20",x"00",x"40",x"C0",x"21",
    x"80",x"20",x"22",x"80",x"20",x"20",x"80",x"00",
    x"00",x"00",x"00",x"63",x"00",x"00",x"20",x"80",
    x"80",x"00",x"A3",x"00",x"E3",x"00",x"00",x"01",
    x"00",x"00",x"00",x"20",x"40",x"24",x"00",x"00",
    x"00",x"00",x"00",x"00",x"40",x"00",x"40",x"00",
    x"00",x"20",x"20",x"00",x"00",x"40",x"00",x"00",
    x"00",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",
    x"A0",x"00",x"00",x"40",x"80",x"00",x"00",x"00",
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",
    x"A0",x"00",x"00",x"40",x"80",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"0C",x"0D",x"0D",x"0E",x"08",x"08",x"08",x"0D",
    x"00",x"E0",x"00",x"00",x"E0",x"00",x"00",x"E0",
    x"00",x"00",x"E0",x"00",x"00",x"E0",x"00",x"00",
    x"E0",x"00",x"44",x"60",x"40",x"A0",x"FF",x"00",
    x"44",x"60",x"40",x"E0",x"00",x"44",x"60",x"00",
    x"60",x"40",x"20",x"FF",x"00",x"80",x"20",x"00",
    x"E0",x"FF",x"00",x"E0",x"00",x"44",x"60",x"40",
    x"A0",x"FF",x"00",x"44",x"60",x"40",x"E0",x"00",
    x"20",x"44",x"60",x"40",x"20",x"40",x"20",x"40",
    x"20",x"40",x"20",x"40",x"40",x"40",x"20",x"40",
    x"40",x"3F",x"40",x"20",x"40",x"3F",x"40",x"E0",
    x"00",x"44",x"60",x"40",x"A0",x"FF",x"00",x"44",
    x"60",x"40",x"60",x"00",x"7F",x"7F",x"44",x"A0",
    x"60",x"40",x"E0",x"FF",x"00",x"44",x"60",x"40",
    x"7F",x"60",x"00",x"00",x"7F",x"40",x"E0",x"00",
    x"BF",x"44",x"00",x"A0",x"E3",x"20",x"A0",x"20",
    x"C0",x"80",x"20",x"FF",x"00",x"00",x"60",x"60",
    x"FF",x"20",x"E0",x"00",x"3C",x"40",x"40",x"20",
    x"00",x"40",x"20",x"00",x"40",x"20",x"00",x"40",
    x"00",x"00",x"00",x"40",x"E0",x"FF",x"3C",x"C0",
    x"20",x"00",x"C0",x"20",x"00",x"C0",x"00",x"C0",
    x"E0",x"00",x"BF",x"40",x"20",x"00",x"3C",x"80",
    x"20",x"00",x"80",x"20",x"00",x"80",x"20",x"00",
    x"80",x"00",x"80",x"00",x"80",x"00",x"E0",x"00",
    x"BF",x"40",x"20",x"00",x"3C",x"80",x"20",x"00",
    x"80",x"20",x"00",x"80",x"20",x"00",x"80",x"00",
    x"44",x"00",x"E0",x"20",x"E0",x"00",x"80",x"C0",
    x"A0",x"FF",x"00",x"00",x"E0",x"FF",x"00",x"00",
    x"A0",x"FF",x"3C",x"80",x"20",x"00",x"80",x"20",
    x"00",x"80",x"00",x"80",x"E0",x"00",x"BF",x"44",
    x"20",x"A0",x"40",x"20",x"40",x"20",x"40",x"20",
    x"40",x"20",x"40",x"40",x"40",x"20",x"40",x"40",
    x"3F",x"40",x"20",x"40",x"00",x"3F",x"A0",x"40",
    x"00",x"00",x"62",x"00",x"60",x"FF",x"00",x"80",
    x"60",x"40",x"E0",x"FF",x"40",x"00",x"3F",x"04",
    x"40",x"60",x"40",x"FF",x"00",x"44",x"00",x"A0",
    x"62",x"00",x"A0",x"80",x"60",x"FF",x"00",x"C0",
    x"60",x"40",x"20",x"FF",x"40",x"44",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"A0",x"E3",x"23",
    x"63",x"E3",x"A3",x"62",x"20",x"60",x"60",x"00",
    x"60",x"FF",x"00",x"00",x"60",x"60",x"00",x"60",
    x"44",x"00",x"A0",x"62",x"00",x"A0",x"80",x"60",
    x"FF",x"00",x"C0",x"60",x"40",x"20",x"FF",x"40",
    x"E0",x"00",x"00",x"60",x"20",x"40",x"04",x"40",
    x"3F",x"00",x"60",x"20",x"60",x"60",x"80",x"00",
    x"60",x"FF",x"00",x"C0",x"A0",x"A0",x"FF",x"60",
    x"00",x"00",x"60",x"00",x"20",x"FF",x"00",x"80",
    x"60",x"40",x"E0",x"FF",x"40",x"00",x"60",x"00",
    x"62",x"40",x"FF",x"00",x"00",x"60",x"00",x"63",
    x"00",x"20",x"FF",x"00",x"80",x"60",x"40",x"E0",
    x"FF",x"40",x"00",x"00",x"60",x"00",x"20",x"FF",
    x"00",x"80",x"60",x"40",x"E0",x"FF",x"40",x"20",
    x"00",x"04",x"FF",x"00",x"FF",x"00",x"C0",x"C0",
    x"FF",x"00",x"00",x"60",x"00",x"20",x"FF",x"00",
    x"80",x"60",x"40",x"E0",x"FF",x"40",x"20",x"00",
    x"04",x"FE",x"00",x"C0",x"C0",x"FF",x"00",x"20",
    x"A0",x"00",x"00",x"C0",x"00",x"60",x"E0",x"FE",
    x"60",x"C0",x"FF",x"00",x"00",x"60",x"00",x"20",
    x"FF",x"00",x"80",x"60",x"40",x"E0",x"FF",x"40",
    x"20",x"00",x"40",x"04",x"40",x"40",x"60",x"20",
    x"00",x"00",x"60",x"20",x"60",x"60",x"80",x"00",
    x"60",x"FF",x"00",x"C0",x"A0",x"A0",x"FF",x"60",
    x"00",x"00",x"60",x"00",x"20",x"FF",x"00",x"80",
    x"60",x"40",x"E0",x"FF",x"40",x"00",x"60",x"00",
    x"63",x"40",x"FF",x"00",x"00",x"00",x"60",x"00",
    x"20",x"FF",x"00",x"80",x"60",x"40",x"E0",x"FF",
    x"40",x"FF",x"00",x"20",x"FF",x"00",x"80",x"60",
    x"40",x"E0",x"FF",x"40",x"FF",x"60",x"00",x"00",
    x"00",x"00",x"20",x"FF",x"00",x"80",x"60",x"40",
    x"E0",x"FF",x"40",x"FF",x"00",x"60",x"FF",x"44",
    x"60",x"40",x"7F",x"60",x"60",x"FF",x"60",x"80",
    x"40",x"00",x"00",x"60",x"FF",x"00",x"00",x"60",
    x"FE",x"60",x"FF",x"00",x"FE",x"00",x"60",x"FF",
    x"00",x"00",x"60",x"FE",x"60",x"FF",x"00",x"FE",
    x"FE",x"00",x"FE",x"20",x"3F",x"BF",x"20",x"FE",
    x"20",x"20",x"20",x"00",x"00",x"00",x"FD",x"60",
    x"C0",x"E0",x"BF",x"40",x"FF",x"00",x"00",x"40",
    x"FD",x"00",x"FD",x"20",x"20",x"FD",x"20",x"7F",
    x"20",x"FD",x"BF",x"C0",x"20",x"20",x"C0",x"00",
    x"00",x"00",x"20",x"00",x"00",x"FD",x"60",x"C0",
    x"E0",x"BF",x"40",x"FF",x"00",x"00",x"40",x"FD",
    x"00",x"FD",x"20",x"FD",x"20",x"20",x"E0",x"FD",
    x"C0",x"E0",x"7F",x"20",x"FD",x"BF",x"C0",x"20",
    x"20",x"C0",x"00",x"00",x"00",x"20",x"00",x"00",
    x"FD",x"60",x"C0",x"E0",x"BF",x"40",x"FF",x"00",
    x"40",x"80",x"00",x"00",x"FD",x"00",x"FE",x"00",
    x"6F",x"61",x"0A",x"00",x"0D",x"00",x"45",x"41",
    x"00",x"00",x"00",x"00",x"54",x"41",x"3A",x"41",
    x"0D",x"00",x"41",x"0D",x"41",x"57",x"45",x"00",
    x"41",x"54",x"0A",x"00",x"53",x"52",x"0A",x"00",
    x"53",x"4B",x"00",x"00",x"00",x"00",x"32",x"36",
    x"41",x"45",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );

  CONSTANT INIT20_3 : type_mem:=(
    x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",
    x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",
    x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"04",x"A0",x"00",x"02",x"00",x"00",x"00",x"00",
    x"80",x"03",x"00",x"80",x"01",x"00",x"80",x"00",
    x"00",x"00",x"04",x"00",x"01",x"0E",x"00",x"00",
    x"00",x"03",x"78",x"03",x"78",x"00",x"00",x"4F",
    x"00",x"00",x"00",x"9E",x"00",x"00",x"60",x"00",
    x"00",x"00",x"00",x"08",x"00",x"08",x"00",x"00",
    x"01",x"01",x"07",x"01",x"00",x"00",x"00",x"00",
    x"00",x"00",x"08",x"10",x"18",x"20",x"28",x"30",
    x"38",x"00",x"13",x"00",x"00",x"00",x"00",x"00",
    x"01",x"07",x"13",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"08",x"10",x"18",x"20",x"28",x"30",
    x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"1E",x"1E",x"1E",x"1E",
    x"9E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",
    x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",
    x"E8",x"40",x"A0",x"1C",x"FC",x"FC",x"FC",x"14",
    x"00",x"08",x"00",x"00",x"08",x"00",x"00",x"08",
    x"00",x"00",x"08",x"00",x"00",x"08",x"00",x"00",
    x"08",x"00",x"00",x"04",x"00",x"04",x"FE",x"00",
    x"00",x"06",x"00",x"08",x"00",x"00",x"06",x"08",
    x"04",x"00",x"04",x"FE",x"00",x"00",x"01",x"00",
    x"00",x"F8",x"00",x"08",x"00",x"00",x"04",x"00",
    x"01",x"FE",x"00",x"00",x"06",x"00",x"08",x"00",
    x"04",x"00",x"04",x"00",x"44",x"00",x"0C",x"00",
    x"0E",x"00",x"0D",x"00",x"00",x"00",x"03",x"00",
    x"00",x"C1",x"00",x"05",x"00",x"EA",x"00",x"08",
    x"00",x"00",x"04",x"00",x"01",x"FE",x"00",x"00",
    x"06",x"00",x"40",x"03",x"D0",x"C9",x"00",x"04",
    x"04",x"00",x"01",x"FE",x"00",x"00",x"06",x"00",
    x"C9",x"40",x"04",x"02",x"D0",x"02",x"08",x"00",
    x"A0",x"00",x"03",x"06",x"58",x"00",x"04",x"1C",
    x"0D",x"00",x"04",x"FE",x"00",x"00",x"01",x"08",
    x"F7",x"04",x"08",x"00",x"00",x"00",x"00",x"50",
    x"02",x"00",x"FF",x"02",x"00",x"40",x"02",x"00",
    x"02",x"02",x"00",x"00",x"80",x"FD",x"00",x"00",
    x"FF",x"02",x"00",x"50",x"02",x"00",x"02",x"00",
    x"08",x"00",x"A0",x"00",x"50",x"01",x"00",x"00",
    x"FF",x"01",x"00",x"60",x"01",x"00",x"D0",x"01",
    x"00",x"01",x"00",x"01",x"00",x"01",x"08",x"00",
    x"A0",x"00",x"50",x"01",x"00",x"00",x"FF",x"01",
    x"00",x"20",x"01",x"00",x"D0",x"01",x"00",x"01",
    x"00",x"01",x"06",x"2D",x"04",x"00",x"00",x"00",
    x"04",x"FE",x"00",x"00",x"80",x"F8",x"00",x"00",
    x"80",x"FE",x"00",x"00",x"FF",x"01",x"00",x"50",
    x"01",x"00",x"01",x"00",x"08",x"00",x"98",x"00",
    x"04",x"04",x"00",x"44",x"00",x"0C",x"00",x"0E",
    x"00",x"0D",x"00",x"00",x"00",x"03",x"00",x"00",
    x"C1",x"00",x"05",x"00",x"01",x"EA",x"06",x"00",
    x"03",x"08",x"C0",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"00",x"FF",x"00",
    x"00",x"04",x"02",x"FD",x"00",x"00",x"03",x"06",
    x"D0",x"08",x"04",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"00",x"01",x"03",
    x"03",x"03",x"03",x"03",x"03",x"00",x"50",x"10",
    x"20",x"40",x"58",x"E8",x"00",x"04",x"06",x"00",
    x"01",x"FE",x"00",x"00",x"5F",x"58",x"14",x"57",
    x"00",x"03",x"06",x"D8",x"08",x"04",x"00",x"04",
    x"FE",x"00",x"00",x"01",x"00",x"00",x"F8",x"00",
    x"08",x"00",x"C3",x"53",x"00",x"00",x"00",x"03",
    x"FF",x"20",x"04",x"00",x"06",x"1C",x"04",x"00",
    x"04",x"FE",x"00",x"00",x"01",x"08",x"F7",x"04",
    x"15",x"08",x"06",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"03",x"06",x"1C",
    x"F0",x"02",x"DD",x"00",x"03",x"06",x"08",x"08",
    x"00",x"04",x"FE",x"00",x"00",x"01",x"00",x"00",
    x"F8",x"00",x"1C",x"1F",x"06",x"00",x"04",x"FE",
    x"00",x"00",x"01",x"00",x"00",x"F8",x"00",x"00",
    x"80",x"00",x"08",x"13",x"1C",x"13",x"18",x"19",
    x"FA",x"1C",x"08",x"06",x"00",x"04",x"FE",x"00",
    x"00",x"01",x"00",x"00",x"F8",x"00",x"00",x"80",
    x"00",x"F1",x"13",x"18",x"19",x"FC",x"00",x"00",
    x"02",x"08",x"00",x"19",x"13",x"10",x"02",x"C5",
    x"10",x"18",x"F9",x"1D",x"08",x"06",x"00",x"04",
    x"FE",x"00",x"00",x"01",x"00",x"00",x"F8",x"00",
    x"00",x"00",x"00",x"00",x"04",x"03",x"10",x"10",
    x"0D",x"20",x"02",x"00",x"06",x"1C",x"04",x"00",
    x"04",x"FE",x"00",x"00",x"01",x"08",x"F7",x"04",
    x"15",x"08",x"06",x"00",x"04",x"FE",x"00",x"00",
    x"01",x"00",x"00",x"F8",x"00",x"03",x"06",x"19",
    x"30",x"02",x"DA",x"00",x"17",x"08",x"06",x"00",
    x"04",x"FE",x"00",x"00",x"01",x"00",x"00",x"F8",
    x"00",x"2E",x"00",x"04",x"FE",x"00",x"00",x"01",
    x"00",x"00",x"F8",x"00",x"23",x"06",x"09",x"1B",
    x"0C",x"00",x"04",x"FE",x"00",x"00",x"01",x"00",
    x"00",x"F8",x"00",x"14",x"00",x"01",x"FE",x"00",
    x"06",x"00",x"D0",x"FF",x"07",x"0A",x"02",x"01",
    x"00",x"00",x"00",x"01",x"FE",x"00",x"00",x"0D",
    x"FF",x"0A",x"F8",x"00",x"FB",x"00",x"01",x"FE",
    x"00",x"00",x"0D",x"F4",x"0A",x"F8",x"00",x"F0",
    x"09",x"00",x"07",x"FF",x"FD",x"FC",x"00",x"02",
    x"FF",x"08",x"FF",x"08",x"06",x"13",x"FB",x"01",
    x"00",x"01",x"FC",x"01",x"FA",x"00",x"43",x"18",
    x"F1",x"00",x"EF",x"FF",x"FF",x"EC",x"08",x"FC",
    x"FF",x"E8",x"FC",x"18",x"FF",x"08",x"00",x"08",
    x"00",x"01",x"00",x"06",x"13",x"DC",x"01",x"00",
    x"01",x"FC",x"01",x"FA",x"00",x"24",x"18",x"D2",
    x"00",x"D0",x"FF",x"CE",x"FF",x"FF",x"08",x"CA",
    x"08",x"08",x"FB",x"FF",x"C5",x"FC",x"18",x"FF",
    x"08",x"00",x"08",x"00",x"01",x"00",x"06",x"13",
    x"B9",x"01",x"00",x"01",x"FC",x"01",x"FA",x"00",
    x"18",x"18",x"02",x"18",x"AD",x"00",x"91",x"00",
    x"74",x"64",x"0D",x"00",x"00",x"00",x"43",x"4D",
    x"00",x"00",x"00",x"00",x"20",x"4E",x"20",x"53",
    x"00",x"00",x"4E",x"00",x"53",x"52",x"0A",x"00",
    x"53",x"45",x"0D",x"00",x"54",x"52",x"0D",x"00",
    x"54",x"0A",x"00",x"00",x"00",x"00",x"33",x"37",
    x"42",x"46",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
    );


  
  SIGNAL wr : unsigned(0 TO 3);
  SIGNAL dr,dw : uv32;

  FUNCTION selvar (
    CONSTANT i5  : type_mem;
    CONSTANT i20 : type_mem) RETURN type_mem IS
  BEGIN
    IF VAR=5 THEN
      RETURN i5;
    ELSE
      RETURN i20;
    END IF;
  END FUNCTION selvar;
  SIGNAL mem0 : type_mem:=selvar(INIT5_0,INIT20_0);
  SIGNAL mem1 : type_mem:=selvar(INIT5_1,INIT20_1);
  SIGNAL mem2 : type_mem:=selvar(INIT5_2,INIT20_2);
  SIGNAL mem3 : type_mem:=selvar(INIT5_3,INIT20_3);
  
  
--------------------------------------------------------------------------------
    
BEGIN

  wr<=mem_w.be WHEN mem_w.req='1' AND mem_w.wr='1' ELSE "0000";

  memproc:PROCESS  (clk)
  BEGIN
    IF rising_edge(clk) THEN
      dr(31 DOWNTO 24)<=mem0(to_integer(mem_w.a(11 DOWNTO 2)));
      IF wr(0)='1' THEN
        mem0(to_integer(mem_w.a(12 DOWNTO 2)))<=dw(31 DOWNTO 24);
      END IF;

      dr(23 DOWNTO 16)<=mem1(to_integer(mem_w.a(11 DOWNTO 2)));
      IF wr(1)='1' THEN
        mem1(to_integer(mem_w.a(12 DOWNTO 2)))<=dw(23 DOWNTO 16);
      END IF;
      
      dr(15 DOWNTO 8)<=mem2(to_integer(mem_w.a(11 DOWNTO 2)));
      IF wr(2)='1' THEN
        mem2(to_integer(mem_w.a(12 DOWNTO 2)))<=dw(15 DOWNTO 8);
      END IF;

      dr(7 DOWNTO 0)<=mem3(to_integer(mem_w.a(11 DOWNTO 2)));
      IF wr(3)='1' THEN
        mem3(to_integer(mem_w.a(12 DOWNTO 2)))<=dw(7 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS memproc;

  mem_r.dr<=dr;
  dw<=mem_w.dw;
  
  mem_r.ack<='1';

END ARCHITECTURE ts;
